module regfile(rd_1, rd_2, rr_1, rr_2, wr, wd, reg_write, clk);
    output reg [31:0] rd_1;
    output reg [31:0] rd_2;
    input [4:0]       rr_1;
    input [4:0]       rr_2;
    input [4:0]       wr;
    input [31:0]      wd;
    input             reg_write;
    input             clk;

    reg [31:0]        reg_file [31:0];
    
    initial begin
        reg_file[00] = 32'b00000000000000000000000000000000;
        reg_file[01] = 32'b00000000000000000000000000000001;
        reg_file[02] = 32'b00000000000000000000000000000010;
        reg_file[03] = 32'b00000000000000000000000000000011;
        reg_file[04] = 32'b00000000000000000000000000000100;
        reg_file[05] = 32'b00000000000000000000000000000101;
        reg_file[06] = 32'b00000000000000000000000000000110;
        reg_file[07] = 32'b00000000000000000000000000000111;
        reg_file[08] = 32'b00000000000000000000000000001000;
        reg_file[09] = 32'b00000000000000000000000000001001;
        reg_file[10] = 32'b00000000000000000000000000001010;
        reg_file[11] = 32'b00000000000000000000000000001011;
        reg_file[12] = 32'b00000000000000000000000000001100;
        reg_file[13] = 32'b00000000000000000000000000001101;
        reg_file[14] = 32'b00000000000000000000000000001110;
        reg_file[15] = 32'b00000000000000000000000000001111;
        reg_file[16] = 32'b00000000000000000000000000010000;
        reg_file[17] = 32'b00000000000000000000000000010001;
        reg_file[18] = 32'b00000000000000000000000000010010;
        reg_file[19] = 32'b00000000000000000000000000010011;
        reg_file[20] = 32'b00000000000000000000000000010100;
        reg_file[21] = 32'b00000000000000000000000000010101;
        reg_file[22] = 32'b00000000000000000000000000010110;
        reg_file[23] = 32'b00000000000000000000000000010111;
        reg_file[24] = 32'b00000000000000000000000000011000;
        reg_file[25] = 32'b00000000000000000000000000011001;
        reg_file[26] = 32'b00000000000000000000000000011010;
        reg_file[27] = 32'b00000000000000000000000000011011;
        reg_file[28] = 32'b00000000000000000000000000011100;
        reg_file[29] = 32'b00000000000000000000000000011101;
        reg_file[30] = 32'b00000000000000000000000000011110;
        reg_file[31] = 32'b00000000000000000000000000011111;

    end
    
    always @ (posedge clk, reg_write) begin
        rd_1 = reg_file[rr_1];
        rd_2 = reg_file[rr_2];
        if (reg_write) begin
            reg_file[wr] = wd;
            // $strobe("(:regfile (:wr %d :wd %d))", wr, wd); 
        end
            
        // $strobe("(:regfile (:rr1 %d :rr2 %d :rd1 %d :rd2 %d))", rr_1, rr_2, rd_1, rd_2);
    end

endmodule