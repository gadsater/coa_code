module not_gate(y, x);
	output y;
	input x;
		
	assign y = ~x;
endmodule
	