module buf_i1(y, x);
	output y;
	input x;
		
	assign y = x;
endmodule
	
