module dummy_tb ();
	string s1;
endmodule
	