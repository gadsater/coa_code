module instr_mem(data, addr, clk);
    output reg [31:0] data;
    input [31:0]      addr;
    input             clk;

    reg [7:0]         mem [127:0];

    initial begin
        mem[000] = 8'b00000000;
        mem[001] = 8'b00000001;
        mem[002] = 8'b11111000;
        mem[003] = 8'b00100000;

        mem[004] = 8'b00000000;
        mem[005] = 8'b00100001;
        mem[006] = 8'b11110000;
        mem[007] = 8'b00100000;

        mem[008] = 8'b00000000;
        mem[009] = 8'b00100010;
        mem[010] = 8'b11101000;
        mem[011] = 8'b00100000;

        mem[012] = 8'b00000000;
        mem[013] = 8'b01000011;
        mem[014] = 8'b11100000;
        mem[015] = 8'b00100000;

        mem[016] = 8'b00000000;
        mem[017] = 8'b01100101;
        mem[018] = 8'b11011000;
        mem[019] = 8'b00100000;

        mem[020] = 8'b00000000;
        mem[021] = 8'b00000000;
        mem[022] = 8'b00000000;
        mem[023] = 8'b00000000;
        mem[024] = 8'b00000000;
        mem[025] = 8'b00000000;
        mem[026] = 8'b00000000;
        mem[027] = 8'b00000000;
        mem[028] = 8'b00000000;
        mem[029] = 8'b00000000;
        mem[030] = 8'b00000000;
        mem[031] = 8'b00000000;
        mem[032] = 8'b00000000;
        mem[033] = 8'b00000000;
        mem[034] = 8'b00000000;
        mem[035] = 8'b00000000;
        mem[036] = 8'b00000000;
        mem[037] = 8'b00000000;
        mem[038] = 8'b00000000;
        mem[039] = 8'b00000000;
        mem[040] = 8'b00000000;
        mem[041] = 8'b00000000;
        mem[042] = 8'b00000000;
        mem[043] = 8'b00000000;
        mem[044] = 8'b00000000;
        mem[045] = 8'b00000000;
        mem[046] = 8'b00000000;
        mem[047] = 8'b00000000;
        mem[048] = 8'b00000000;
        mem[049] = 8'b00000000;
        mem[050] = 8'b00000000;
        mem[051] = 8'b00000000;
        mem[052] = 8'b00000000;
        mem[053] = 8'b00000000;
        mem[054] = 8'b00000000;
        mem[055] = 8'b00000000;
        mem[056] = 8'b00000000;
        mem[057] = 8'b00000000;
        mem[058] = 8'b00000000;
        mem[059] = 8'b00000000;
        mem[060] = 8'b00000000;
        mem[061] = 8'b00000000;
        mem[062] = 8'b00000000;
        mem[063] = 8'b00000000;
        mem[064] = 8'b00000000;
        mem[065] = 8'b00000000;
        mem[066] = 8'b00000000;
        mem[067] = 8'b00000000;
        mem[068] = 8'b00000000;
        mem[069] = 8'b00000000;
        mem[070] = 8'b00000000;
        mem[071] = 8'b00000000;
        mem[072] = 8'b00000000;
        mem[073] = 8'b00000000;
        mem[074] = 8'b00000000;
        mem[075] = 8'b00000000;
        mem[076] = 8'b00000000;
        mem[077] = 8'b00000000;
        mem[078] = 8'b00000000;
        mem[079] = 8'b00000000;
        mem[080] = 8'b00000000;
        mem[081] = 8'b00000000;
        mem[082] = 8'b00000000;
        mem[083] = 8'b00000000;
        mem[084] = 8'b00000000;
        mem[085] = 8'b00000000;
        mem[086] = 8'b00000000;
        mem[087] = 8'b00000000;
        mem[088] = 8'b00000000;
        mem[089] = 8'b00000000;
        mem[090] = 8'b00000000;
        mem[091] = 8'b00000000;
        mem[092] = 8'b00000000;
        mem[093] = 8'b00000000;
        mem[094] = 8'b00000000;
        mem[095] = 8'b00000000;
        mem[096] = 8'b00000000;
        mem[097] = 8'b00000000;
        mem[098] = 8'b00000000;
        mem[099] = 8'b00000000;
        mem[100] = 8'b00000000;
        mem[101] = 8'b00000000;
        mem[102] = 8'b00000000;
        mem[103] = 8'b00000000;
        mem[104] = 8'b00000000;
        mem[105] = 8'b00000000;
        mem[106] = 8'b00000000;
        mem[107] = 8'b00000000;
        mem[108] = 8'b00000000;
        mem[109] = 8'b00000000;
        mem[110] = 8'b00000000;
        mem[111] = 8'b00000000;
        mem[112] = 8'b00000000;
        mem[113] = 8'b00000000;
        mem[114] = 8'b00000000;
        mem[115] = 8'b00000000;
        mem[116] = 8'b00000000;
        mem[117] = 8'b00000000;
        mem[118] = 8'b00000000;
        mem[119] = 8'b00000000;
        mem[120] = 8'b00000000;
        mem[121] = 8'b00000000;
        mem[122] = 8'b00000000;
        mem[123] = 8'b00000000;
        mem[124] = 8'b00000000;
        mem[125] = 8'b00000000;
        mem[126] = 8'b00000000;
        mem[127] = 8'b00000000;
    end
    always @ (posedge clk) begin
       data = {mem[addr[6:0] + 7'b0000000], 
               mem[addr[6:0] + 7'b0000001],
               mem[addr[6:0] + 7'b0000010],
               mem[addr[6:0] + 7'b0000011]};
        // $strobe("(:instr-mem (:addr %d :data %d))", addr, data); 

    end
endmodule